library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity InstructionMemory is
    Port ( Address : in  STD_LOGIC_VECTOR (5 downto 0);
           rst : in  STD_LOGIC;
           Instruction : out  STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture syn of InstructionMemory is

type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);                 
signal ROM : rom_type:= ("00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000","00000001000000000000000000000000",
								 "00000001000000000000000000000000",
								 "10010000000100000000000000010000",
								 "10110010000100000010000000000110","01111111111111111111111111110100",
								 "10100010000100000000000000010010","00010000101111111111111111111000",--"10000001110000000010000000000100",
								 "10100100000001000110000000000001","10100000000100000000000000010010",
								 "10100100000001000000000000011000",
								 "00000001000000000000000000000000","10000001110000111110000000000010",
								 "00000001000000000000000000000000","00101100100000000000000000000100",
								 "10000000101001000100000000011001","10100010000100000010000000000000",
								 "10100000000100000010000000000000","10110000000100000010000000001100",
								 "01000000000000000000000000001110");
								 --"00000000000000000000000000000000","10011110000001000100000000010000",
								 --"10101110100001010100000000010110","10101101001011010011000000010100",--"10101100100001010100000000010101",								
								 --"10101011001011010011000000010011","10101000000100000010111111111111",
								 --"10100110100101000000000000010001","10100110100010000010011110101000",
								 --"10010000001001000100000000010010","10100100000001000010000000010000",
								 --"10100010000100000010000000010001","10100000000100000010000000001111");                        

begin

process(rst,Address,ROM)

begin

if rst='1' then
	Instruction<=(others=>'0');
else
	Instruction<=ROM(conv_integer(Address));
end if;

end process;

end syn;