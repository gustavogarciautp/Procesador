library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

entity InstructionMemory is
    Port ( Address : in  STD_LOGIC_VECTOR (5 downto 0);
           rst : in  STD_LOGIC;
           Instruction : out  STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory;

architecture syn of InstructionMemory is

type rom_type is array (63 downto 0) of std_logic_vector (31 downto 0);                 
signal ROM : rom_type:= ("00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",
								 "00000000000000000000000000000000","00000000000000000000000000000000",								
								 "00000000000000000000000000000000","10011000001000000100000000000010",
								 "10010110001110000100000000000010","10010100001010000100000000000010",
								 "10010010000110000100000000000010","10010000000000000100000000000010",
								 "10000100000100000011111111111001","10000010000100000010000000001000");                          

begin

process(rst,Address,ROM)

begin

if rst='1' then
	Instruction<=(others=>'0');
else
	Instruction<=ROM(conv_integer(Address));
end if;

end process;

end syn;
